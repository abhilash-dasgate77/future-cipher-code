`timescale 1ns / 1ps

module mux_sbmx_sb(a,b,s);
	input [0:15]a,s;
	output [0:15]b;
	assign b[0] = 
endmodule
