`timescale 1ns / 1ps

module or_1bit(
    input a,
    input b,
    output c
    );
	assign c = a | b;
endmodule
